module mips_rom(
    input [31:0] address,
    output reg [31:0] data
);

always @(address) begin
    case(address)
    //Program 1:
    //This sequence of instructions is a LD R2,M[R1+127] (0+127 / 4) = M[31]
     //a LD R3,M[R1+128] (0+128 / 4) = M[32]
     //and an ADD R4,R2,R3 (R4 = R2 + R3)
		/*
     32'h0000_0000: data = 32'b1000_1100_0010_0010_0000_0000_0111_1111;
     32'h0000_0001: data = 32'b1000_1100_0010_0011_0000_0000_1000_0010;
     32'h0000_0002: data= 32'b0000_0000_0100_0011_0010_0000_0010_0000;
     32'h0000_001F: data = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
     32'h0000_0020: data = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
	*/
    /*32'h0000_0000: data = 32'b1000_1100_0000_0001_0000_0000_0111_1111; //LD R1,M[31]
    32'h0000_0001: data = 32'b1000_1100_0000_0010_0000_0000_1000_0010; //LD R2,M[32]
    32'h0000_0002: data = 32'b0000_0000_0010_0010_0000_1000_0010_0010; //SUB R1,R1,R2
    32'h0000_0003: data = 32'b0001_0000_0000_0001_0000_0000_0000_0001; //BEQ R0,R1, DONE
    32'h0000_0004: data = 32'b0000_1000_0000_0000_0000_0000_0000_0010; //JMP, 0x0008
    32'h0000_0005: data = 32'b0000_1000_0000_0000_0000_0000_0000_0101; //JMP, 0x0005 (INF. LOOP)
    32'h0000_001F: data = 32'b0000_0000_0000_0000_0000_0000_0000_0101;
    32'h0000_0020: data = 32'b0000_0000_0000_0000_0000_0000_0000_0001;    
*/
	 32'h0000_0000: data = 32'b1000_1100_0000_0001_0000_0000_0111_1111; //LD R1,M[31]
	 32'h0000_0001: data = 32'b1000_1100_0000_0010_0000_0000_1000_0010; //LD R2,M[32]
	 32'h0000_0002: data = 32'b1000_1100_0000_0011_0000_0000_1000_0100; //LD R3,M[33]
	 32'h0000_0003: data = 32'b1000_1100_0000_0100_0000_0000_1000_1000; //LD R4,M[34]
	 32'h0000_0004: data = 32'b1000_1100_0000_0101_0000_0000_1000_1100; //LD R5,M[35]
	 32'h0000_0005: data = 32'b1010_1100_0010_0011_0000_0000_0000_0000; //SW M[DESLSB],R3
	 32'h0000_0006: data = 32'b1010_1100_0010_0010_0000_0000_0001_0000; //SW M[DESMSB],R2
	 32'h0000_0007: data = 32'b1010_1100_0010_0100_0000_0000_0010_0000; //SW M[KEYLSB],R4
	 32'h0000_0008: data = 32'b1010_1100_0010_0101_0000_0000_0011_0000; //SW M[KEYMSB],R5
	 32'h0000_001F: data = 32'b00000000000000110000100000000000; 		  //M[31]
	 32'h0000_0020: data = 32'b10001001101010111100110111101111; 		  //M[32]
	 32'h0000_0021: data = 32'b00000001001000110100010101100111; 		  //M[33]
	 32'h0000_0022: data = 32'h13345779; 									     //M[34]
	 32'h0000_0023: data = 32'h9BBCDFF1; 										  //M[35]




    default: data = 32'hFFFF_FFFF;
    endcase
end


endmodule
